library verilog;
use verilog.vl_types.all;
entity DataOut_v1_vlg_vec_tst is
end DataOut_v1_vlg_vec_tst;
