library verilog;
use verilog.vl_types.all;
entity Alu_v1_vlg_vec_tst is
end Alu_v1_vlg_vec_tst;
