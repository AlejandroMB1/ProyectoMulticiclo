library verilog;
use verilog.vl_types.all;
entity MuxPc_v1_vlg_vec_tst is
end MuxPc_v1_vlg_vec_tst;
