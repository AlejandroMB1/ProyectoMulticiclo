library verilog;
use verilog.vl_types.all;
entity PC_v1_vlg_vec_tst is
end PC_v1_vlg_vec_tst;
