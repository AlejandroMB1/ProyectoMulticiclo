library verilog;
use verilog.vl_types.all;
entity Arquitectura_v1_vlg_vec_tst is
end Arquitectura_v1_vlg_vec_tst;
