library verilog;
use verilog.vl_types.all;
entity IR_v1_vlg_vec_tst is
end IR_v1_vlg_vec_tst;
